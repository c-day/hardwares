
module MEM(PCSrc, readData, memRead, memWrite, sawBranch, branchOp, clk, writeData, address);
  input [15:0] writeData;
  input sawBranch, memRead, memWrite, clk;
  input [2:0] branchOp;
  output [15:0] readData;
  output PCSrc;
  inout [15:0] address;
  
  DM dataMem(.clk(clk),.addr(address),.re(memRead),.we(memWrite),.wrt_data(writeData),.rd_data(readData));
  
  branchLogic branchLogic(.PCSrc(PCSrc), .takeBranch(sawBranch), .branchOp(branchOp));
  
  
endmodule