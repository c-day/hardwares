/*******************************************************************************
* ECE 552 ALU
* Author: Craig Day and Ethan Massey
*
* The ALU accepts 2 16 bit sources (src0, src1) and will perform the operation
* specified by the 4 bit control signal (ctrl).  It will return the result on 
* a 16 bit bus (dst) and set overflow (ov) and zero (zr) flags accordingly. When
* a shit is to be performed, src0 will be shifted by an amount specified in the
* shamt parameter.
*
* Parameters:
* src0 - input used for all operations
* src1 - input used in any two-op operations
* ctrl - the control signal specifying the operation to be performed
* shamt - the amount to shift by if a shift is being performed
* 
* Returns:
* dst - the result of the operation specified by ctrl
* ov - contains 1 on overflow, 0 otherwise
* zr - contains 1 if result is 0, 0 otherwise
*******************************************************************************/

module ALU(dst, ov, zr, src0, src1, ctrl, shamt);
	input [15:0] src0, src1;
	input [3:0] ctrl;
	input [3:0] shamt;
	output [15:0] dst;
	output ov, zr;

	// Use parameters so that the opcodes can be specified by higher
	// level modules.  
	parameter addOp = 3'b000;
	parameter subOp = 3'b001;
	parameter andOp = 3'b010;
	parameter norOp = 3'b011;
	parameter sllOp = 3'b100;
	parameter srlOp = 3'b101;
	parameter sraOp = 3'b110;
	parameter lhbOp = 3'b111;

	//signed wire to contain the right arithmatic shift value	
	wire signed [15:0] sra;
	
	// do the right arathmatic shift using the signed bus,
	// forces the MSB to behave correctly
	assign sra = src0 >>> shamt;
	
	//parallel_case
	assign 	{ov, dst} = (ctrl == addOp) ? src0 + src1 :
											(ctrl == subOp) ? src0 - src1 :
											(ctrl == andOp) ? {1'b0, src0 & src1} :
											(ctrl == norOp) ? {1'b0, ~(src0 | src1)} :
											(ctrl == sllOp) ? {1'b0, src0 << shamt} :
											(ctrl == srlOp) ? {1'b0, src0 >> shamt} :
											(ctrl == sraOp) ? {1'b0, sra} :	
											(ctrl == lhbOp) ? {1'b0, {src0[15:8], 8'd0} | src1} :
											17'd0;
	
// nor all of the bits together, will set zr to 1 only when all bits of result are 0
	assign zr = ~|dst;

endmodule